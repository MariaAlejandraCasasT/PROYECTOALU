library verilog;
use verilog.vl_types.all;
entity ALU_P_vlg_vec_tst is
end ALU_P_vlg_vec_tst;
