library verilog;
use verilog.vl_types.all;
entity ALUFull_P_vlg_vec_tst is
end ALUFull_P_vlg_vec_tst;
